library ieee;
use ieee.std_logic_1164.all;

use work.types.all;

entity SGMII_SI_data is
  
  port (
    entry : in  integer;
    addr  : out slv_12_t;
    data  : out slv_8_t);

end entity SGMII_SI_data;

architecture behavioral of SGMII_SI_data is

  --Upper 12  bits are addr, lower 12 are data
  constant writes : slv20_array_t(0 to 464) := (x"B24C0",
                                              x"B2500",
                                              x"54001",
                                              x"00600",
                                              x"00700",
                                              x"00800",
                                              x"00B68",
                                              x"01602",
                                              x"017DC",
                                              x"018EE",
                                              x"019DD",
                                              x"01ADF",
                                              x"02B02",
                                              x"02C01",
                                              x"02D01",
                                              x"02E38",
                                              x"02F00",
                                              x"03000",
                                              x"03100",
                                              x"03200",
                                              x"03300",
                                              x"03400",
                                              x"03500",
                                              x"03638",
                                              x"03700",
                                              x"03800",
                                              x"03900",
                                              x"03A00",
                                              x"03B00",
                                              x"03C00",
                                              x"03D00",
                                              x"03F11",
                                              x"04004",
                                              x"0410D",
                                              x"04200",
                                              x"04300",
                                              x"04400",
                                              x"0450C",
                                              x"04632",
                                              x"04700",
                                              x"04800",
                                              x"04900",
                                              x"04A32",
                                              x"04B00",
                                              x"04C00",
                                              x"04D00",
                                              x"04E05",
                                              x"04F00",
                                              x"0500F",
                                              x"05103",
                                              x"05200",
                                              x"05300",
                                              x"05400",
                                              x"05503",
                                              x"05600",
                                              x"05700",
                                              x"05800",
                                              x"05901",
                                              x"05AAA",
                                              x"05BAA",
                                              x"05C0A",
                                              x"05D01",
                                              x"05E00",
                                              x"05F00",
                                              x"06000",
                                              x"06100",
                                              x"06200",
                                              x"06300",
                                              x"06400",
                                              x"06500",
                                              x"06600",
                                              x"06700",
                                              x"06800",
                                              x"06900",
                                              x"09202",
                                              x"093A0",
                                              x"09500",
                                              x"09680",
                                              x"09860",
                                              x"09A02",
                                              x"09B60",
                                              x"09D08",
                                              x"09E40",
                                              x"0A020",
                                              x"0A200",
                                              x"0A9A7",
                                              x"0AA61",
                                              x"0AB00",
                                              x"0AC00",
                                              x"0E521",
                                              x"0EA0A",
                                              x"0EB60",
                                              x"0EC00",
                                              x"0ED00",
                                              x"10201",
                                              x"11202",
                                              x"11309",
                                              x"11433",
                                              x"11508",
                                              x"11702",
                                              x"11809",
                                              x"11933",
                                              x"11A08",
                                              x"12602",
                                              x"12709",
                                              x"12833",
                                              x"12909",
                                              x"12B02",
                                              x"12C09",
                                              x"12D33",
                                              x"12E0A",
                                              x"13F00",
                                              x"14000",
                                              x"14140",
                                              x"142FF",
                                              x"20600",
                                              x"20832",
                                              x"20900",
                                              x"20A00",
                                              x"20B00",
                                              x"20C00",
                                              x"20D00",
                                              x"20E01",
                                              x"20F00",
                                              x"21000",
                                              x"21100",
                                              x"21200",
                                              x"21300",
                                              x"21400",
                                              x"21500",
                                              x"21600",
                                              x"21700",
                                              x"21800",
                                              x"21900",
                                              x"21A00",
                                              x"21B00",
                                              x"21C00",
                                              x"21D00",
                                              x"21E00",
                                              x"21F00",
                                              x"22000",
                                              x"22100",
                                              x"22200",
                                              x"22300",
                                              x"22400",
                                              x"22500",
                                              x"22600",
                                              x"22700",
                                              x"22800",
                                              x"22900",
                                              x"22A00",
                                              x"22B00",
                                              x"22C00",
                                              x"22D00",
                                              x"22E00",
                                              x"22F00",
                                              x"2310B",
                                              x"2320B",
                                              x"2330B",
                                              x"2340B",
                                              x"23500",
                                              x"23600",
                                              x"23700",
                                              x"238C0",
                                              x"239DA",
                                              x"23A00",
                                              x"23B00",
                                              x"23C00",
                                              x"23D00",
                                              x"23EC0",
                                              x"25003",
                                              x"25100",
                                              x"25200",
                                              x"25304",
                                              x"25400",
                                              x"25500",
                                              x"25C02",
                                              x"25D00",
                                              x"25E00",
                                              x"25F02",
                                              x"26000",
                                              x"26100",
                                              x"26B41",
                                              x"26C50",
                                              x"26D4F",
                                              x"26E4C",
                                              x"26F4C",
                                              x"2704F",
                                              x"27153",
                                              x"2724D",
                                              x"28A00",
                                              x"28B00",
                                              x"28C00",
                                              x"28D00",
                                              x"28E00",
                                              x"28F00",
                                              x"29000",
                                              x"29100",
                                              x"294B0",
                                              x"29602",
                                              x"29702",
                                              x"29902",
                                              x"29DFA",
                                              x"29E01",
                                              x"29F00",
                                              x"2A9CC",
                                              x"2AA04",
                                              x"2AB00",
                                              x"2B7FF",
                                              x"30200",
                                              x"30300",
                                              x"30400",
                                              x"30500",
                                              x"30607",
                                              x"30700",
                                              x"30800",
                                              x"30900",
                                              x"30A00",
                                              x"30B80",
                                              x"30C00",
                                              x"30D00",
                                              x"30E00",
                                              x"30FEC",
                                              x"31060",
                                              x"31121",
                                              x"31200",
                                              x"31300",
                                              x"314B8",
                                              x"315C6",
                                              x"31692",
                                              x"31700",
                                              x"31800",
                                              x"319C0",
                                              x"31A49",
                                              x"31B6E",
                                              x"31C0A",
                                              x"31D00",
                                              x"31E00",
                                              x"31F8B",
                                              x"32077",
                                              x"321B7",
                                              x"32200",
                                              x"32300",
                                              x"32400",
                                              x"32500",
                                              x"32600",
                                              x"32700",
                                              x"32800",
                                              x"32900",
                                              x"32A00",
                                              x"32B00",
                                              x"32C00",
                                              x"32D00",
                                              x"33800",
                                              x"3391F",
                                              x"33B00",
                                              x"33C00",
                                              x"33D00",
                                              x"33E00",
                                              x"33F00",
                                              x"34000",
                                              x"34100",
                                              x"34200",
                                              x"34300",
                                              x"34400",
                                              x"34500",
                                              x"34600",
                                              x"34700",
                                              x"34800",
                                              x"34900",
                                              x"34A00",
                                              x"34B00",
                                              x"34C00",
                                              x"34D00",
                                              x"34E00",
                                              x"34F00",
                                              x"35000",
                                              x"35100",
                                              x"35200",
                                              x"35900",
                                              x"35A00",
                                              x"35B00",
                                              x"35C00",
                                              x"35D00",
                                              x"35E00",
                                              x"35F00",
                                              x"36000",
                                              x"48700",
                                              x"50813",
                                              x"50922",
                                              x"50A0C",
                                              x"50B0B",
                                              x"50C07",
                                              x"50D3F",
                                              x"50E16",
                                              x"50F2A",
                                              x"51009",
                                              x"51108",
                                              x"51207",
                                              x"5133F",
                                              x"51500",
                                              x"51600",
                                              x"51700",
                                              x"51800",
                                              x"519BC",
                                              x"51A02",
                                              x"51B00",
                                              x"51C00",
                                              x"51D00",
                                              x"51E00",
                                              x"51F80",
                                              x"5212B",
                                              x"52A01",
                                              x"52B01",
                                              x"52C87",
                                              x"52D03",
                                              x"52E19",
                                              x"52F19",
                                              x"53100",
                                              x"53242",
                                              x"53303",
                                              x"53400",
                                              x"53500",
                                              x"53604",
                                              x"53700",
                                              x"53800",
                                              x"53900",
                                              x"53A02",
                                              x"53B03",
                                              x"53C00",
                                              x"53D11",
                                              x"53E06",
                                              x"5890D",
                                              x"58A00",
                                              x"59BFA",
                                              x"59D13",
                                              x"59E24",
                                              x"59F0C",
                                              x"5A00B",
                                              x"5A107",
                                              x"5A23F",
                                              x"5A603",
                                              x"80235",
                                              x"80305",
                                              x"80400",
                                              x"80500",
                                              x"80600",
                                              x"80700",
                                              x"80800",
                                              x"80900",
                                              x"80A00",
                                              x"80B00",
                                              x"80C00",
                                              x"80D00",
                                              x"80E00",
                                              x"80F00",
                                              x"81000",
                                              x"81100",
                                              x"81200",
                                              x"81300",
                                              x"81400",
                                              x"81500",
                                              x"81600",
                                              x"81700",
                                              x"81800",
                                              x"81900",
                                              x"81A00",
                                              x"81B00",
                                              x"81C00",
                                              x"81D00",
                                              x"81E00",
                                              x"81F00",
                                              x"82000",
                                              x"82100",
                                              x"82200",
                                              x"82300",
                                              x"82400",
                                              x"82500",
                                              x"82600",
                                              x"82700",
                                              x"82800",
                                              x"82900",
                                              x"82A00",
                                              x"82B00",
                                              x"82C00",
                                              x"82D00",
                                              x"82E00",
                                              x"82F00",
                                              x"83000",
                                              x"83100",
                                              x"83200",
                                              x"83300",
                                              x"83400",
                                              x"83500",
                                              x"83600",
                                              x"83700",
                                              x"83800",
                                              x"83900",
                                              x"83A00",
                                              x"83B00",
                                              x"83C00",
                                              x"83D00",
                                              x"83E00",
                                              x"83F00",
                                              x"84000",
                                              x"84100",
                                              x"84200",
                                              x"84300",
                                              x"84400",
                                              x"84500",
                                              x"84600",
                                              x"84700",
                                              x"84800",
                                              x"84900",
                                              x"84A00",
                                              x"84B00",
                                              x"84C00",
                                              x"84D00",
                                              x"84E00",
                                              x"84F00",
                                              x"85000",
                                              x"85100",
                                              x"85200",
                                              x"85300",
                                              x"85400",
                                              x"85500",
                                              x"85600",
                                              x"85700",
                                              x"85800",
                                              x"85900",
                                              x"85A00",
                                              x"85B00",
                                              x"85C00",
                                              x"85D00",
                                              x"85E00",
                                              x"85F00",
                                              x"86000",
                                              x"86100",
                                              x"90E02",
                                              x"94300",
                                              x"94901",
                                              x"94A01",
                                              x"94E49",
                                              x"94F02",
                                              x"95E00",
                                              x"A0200",
                                              x"A0307",
                                              x"A0401",
                                              x"A0507",
                                              x"A1400",
                                              x"A1A00",
                                              x"A2000",
                                              x"A2600",
                                              x"B442F",
                                              x"B4600",
                                              x"B470E",
                                              x"B480E",
                                              x"B4A08",
                                              x"B570E",
                                              x"B5801",
                                              x"51401",
                                              x"01C01",
                                              x"54000",
                                              x"B24C3",
                                              x"B2502"
                                              );
begin  -- architecture behavioral

  addr <= writes(entry)(19 downto 8);
  data <= writes(entry)( 7 downto 0);

end architecture behavioral;
